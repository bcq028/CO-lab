`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/10/23 15:21:30
// Design Name: 
// Module Name: controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module controller(
	input wire clk,rst,
	//decode stage
	input wire[5:0] opD,functD,
	output wire pcsrcD,branchD,equalD,jumpD,
	
	//execute stage
	input wire flushE,
	output wire memtoregE,
	output wire[1:0] alusrcE,
	output wire regdstE,regwriteE,	
	output wire[4:0] alucontrolE,

	//mem stage
	output wire memtoregM,memwriteM,
				regwriteM,
	//write back stage
	output wire memtoregW,regwriteW

    );
	
	//decode stage
	wire[3:0] aluopD;
	wire memtoregD,memwriteD,
		regdstD,regwriteD;
	wire [1:0] alusrcD;
	wire[4:0] alucontrolD;

	//execute stage
	wire memwriteE;

	maindec md(
		.op(opD),
		.regwrite(regwriteD),
		.regdst(regdstD),
		.alusrc(alusrcD),
		.branch(branchD),
		.memwrite(memwriteD),
		.memtoreg(memtoregD),
		.jump(jumpD),
		.aluop(aluopD)
    );

	aludec aludec (
		.funct 		(functD		),
		.aluop 		(aluopD		),
		.alucontrol	(alucontrolD)
	);

	assign pcsrcD = branchD & equalD;

	//pipeline registers
	floprc #(11) regE(
		clk,
		rst,
		flushE,
		{memtoregD,memwriteD,alusrcD,regdstD,regwriteD,alucontrolD},
		{memtoregE,memwriteE,alusrcE,regdstE,regwriteE,alucontrolE}
		);
	flopr #(11) regM(
		clk,rst,
		{memtoregE,memwriteE,regwriteE},
		{memtoregM,memwriteM,regwriteM}
		);
	flopr #(11) regW(
		clk,rst,
		{memtoregM,regwriteM},
		{memtoregW,regwriteW}
		);
endmodule
